** Profile: "SCHEMATIC1-control"  [ C:\ORCAD\ORCAD_10.3\proyecto\motor-pspicefiles\schematic1\control.sim ] 

** Creating circuit file "control.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\ORCAD\ORCAD_10.3\proyecto\motor-pspicefiles\schematic1\control\control_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_10.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1s 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
